

class src_seqr extends uvm_sequencer #(trans);

	`uvm_component_utils(src_seqr)
	function new(string name="src_seqr",uvm_component parent);
		super.new(name,parent);
	endfunction


endclass

