

class router_virtual_seqs extends uvm_sequence #(uvm_sequence_item);
	`uvm_object_utils(router_virtual_seqs)  
	
	function new(string name ="router_virtual_seqs");
		super.new(name);
	endfunction
endclass

